package spi_test_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "m_xtn.sv"
`include "s_xtn.sv"

`include "m_agt_cfg.sv"
`include "s_agt_cfg.sv"
`include "spi_env_cfg.sv"

`include "m_drv.sv"
`include "m_mon.sv"
`include "m_seqr.sv"
`include "m_agt.sv"
`include "m_agt_top.sv"
`include "m_seq.sv"

`include "s_drv.sv"
`include "s_mon.sv"
`include "s_seqr.sv"
`include "s_agt.sv"
`include "s_agt_top.sv"
`include "s_seq.sv"

`include "spi_vseqr.sv"
`include "spi_vseqs.sv"
`include "spi_sb.sv"
`include "spi_env.sv"
`include "spi_test.sv"

endpackage