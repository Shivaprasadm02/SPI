class m_seqr extends uvm_sequencer#(m_xtn);

`uvm_component_utils(m_seqr)

function new(string name="m_seqr",uvm_component parent);
	super.new(name,parent);
endfunction 

endclass