class
endclass
